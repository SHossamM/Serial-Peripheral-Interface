library verilog;
use verilog.vl_types.all;
entity Master_tb is
end Master_tb;
